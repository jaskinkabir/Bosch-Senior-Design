PLC_Diag_One_PSU

.TRAN 1ms 100ms
* .AC DEC 100 100 1MEG
.END
